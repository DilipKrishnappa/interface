//module : interface
//static component
interface intf();
  //Declare the signals
  logic [3:0]a,b;
  logic [6:0]y;
endinterface
//end module: interface 
